library verilog;
use verilog.vl_types.all;
entity test_stepmot is
end test_stepmot;
