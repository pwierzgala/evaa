/*****************************************************************************************************************
* Test Bench for Step Motor Controller
* December 2006
*****************************************************************************************************************/


module test_stepmot;
 
 /* Applied test stimuli, corresponding to: reset,mode,	dir, move, phaseout. */

 reg [3:0] test_vec;   
 reg oscena;

 wire [3:0] test_phase;             //output generated by the controller module.
 wire osc,clk_t,clk1;

 integer t;
  
 initial
  begin
     oscena=1'b1;
     t=0;
  end

/* Mapping the test bench varialbles into the main module variables.*/
 stepmot s1_t(                        
         .reset (test_vec[3]),
         .mode (test_vec[2]),
         .dir (test_vec[1]),
         .move (test_vec[0]),
         .phaseout(test_phase)); 
 ufmclk  ufm1(                     //Instantiation  of ufmclk module.
        .oscena (oscena),
        .osc  (osc));
                     
 divider1 d1_t( 
        .osc  (osc),               //Instantiation  of clk divider module.
        .clk  (clk_t),
        .clk1  (clk1));
        
  initial
  
       $monitor("Simulation period:%d,       Test vector:%b,        Test phase:%b",$time,test_vec,test_phase);
        
/* Providing all valid inputs to the main module of Stepper motor */        
always @( negedge clk_t)
     begin
       if(t==0)
            test_vec=4'b0011;       
       if(t==1)
            test_vec=4'b1011;
       if(t==2) 
            test_vec=4'b1011;
       if(t==3)
            test_vec=4'b1011;
       if(t==4)
            test_vec=4'b1011; 
       if(t==5)  
            test_vec=4'b1011;
       if(t==6)
            test_vec=4'b1011;
       if(t==7)
            test_vec=4'b1011;
       if(t==8)
            test_vec=4'b1011;
       if(t==9)
            test_vec=4'b1001;
       if(t==10)
            test_vec=4'b1001;
       if(t==11)
            test_vec=4'b1001;
       if(t==12)
            test_vec=4'b1001;
       if(t==13)
            test_vec=4'b1001;
       if(t==14)
            test_vec=4'b1001;
       if(t==15)
            test_vec=4'b1001;
       if(t==16)
            test_vec=4'b1001;
       if(t==17)
            test_vec=4'b1111;
       if(t==18)
            test_vec=4'b1110;
       if(t==19)
            test_vec=4'b1111;
       if(t==20)
            test_vec=4'b1110;
       if(t==21)
            test_vec=4'b1111;
       if(t==22)
            test_vec=4'b1110;
       if(t==23)
            test_vec=4'b1111;
       if(t==24)
            test_vec=4'b1110;
       if(t==25)
            test_vec=4'b1111;
       if(t==26)
            test_vec=4'b1110;
       if(t==27)
            test_vec=4'b1111;
       if(t==28)
            test_vec=4'b1110;
       if(t==29)
            test_vec=4'b1111;
       if(t==30)
            test_vec=4'b1110;
       if(t==31)
            test_vec=4'b1111;
       if(t==32)
            test_vec=4'b1110;
       if(t==33)
            test_vec=4'b1111;
       if(t==34)
            test_vec=4'b1110;
       if(t==35)
            test_vec=4'b1101;
       if(t==36)
            test_vec=4'b1100;
       if(t==37)
            test_vec=4'b1101;
       if(t==38)
            test_vec=4'b1100;
       if(t==39)
            test_vec=4'b1101;
       if(t==40)
            test_vec=4'b1100;
       if(t==41)
            test_vec=4'b1101;
       if(t==42)
            test_vec=4'b1100;
       if(t==43)
            test_vec=4'b1101;
       if(t==44)
            test_vec=4'b1100;
       if(t==45)
            test_vec=4'b1101;
       if(t==46)
            test_vec=4'b1100;
       if(t==47)
            test_vec=4'b1101;
       if(t==48)
            test_vec=4'b1100;
       if(t==49)
            test_vec=4'b1101;
       if(t==50)
            test_vec=4'b1100;
       if(t==51)
            test_vec=4'b1101;
       if(t==52)
            test_vec=4'b1100;
       if(t==53)
            test_vec=4'b1101;               
                                         
       t=t+1;
    end 
         
/* Process to check the outputs for the corresponding inputs */
always @( posedge clk1) begin
   if (clk_t==1'b1)begin
       
       if(t==1) begin
           if(test_phase== 4'b0111)
           $display ("Output Verified");
           else begin 
           $display ("Error"); 
           $stop;end
           end
                 
       if(t==2) begin
           if(test_phase== 4'b0011)
           $display ("Output Verified");
           else begin 
           $display ("Error"); 
           $stop;end
           end
          
       if(t==3) begin
           if(test_phase== 4'b1011)
           $display ("Output Verified");
           else begin 
           $display ("Error"); 
           $stop; end
           end
                 
       if(t==4) begin
           if(test_phase== 4'b1001)
           $display ("Output Verified");
           else begin
           $display ("Error");
           $stop; end
           end
                 
       if(t==5) begin
           if(test_phase== 4'b1101)
           $display ("Output Verified");
           else begin
           $display ("Error");
           $stop; end
           end
                 
       if(t==6) begin
           if(test_phase== 4'b1100)
           $display ("Output Verified");
           else begin 
           $display ("Error"); 
           $stop; end
           end
              
       if(t==7) begin
           if(test_phase== 4'b1110)
           $display ("Output Verified");
           else begin 
           $display ("Error");
           $stop; end
           end
               
       if(t==8) begin
           if(test_phase== 4'b0110)
           $display ("Output Verified");
           else begin
           $display ("Error");
           $stop; end
           end
    
       if(t==9) begin
           if(test_phase== 4'b0111)
           $display ("Output Verified");
           else begin
           $display ("Error"); 
           $stop; end
           end
   
       if(t==10) begin
           if(test_phase== 4'b0110)
           $display ("Output Verified");
           else begin 
           $display ("Error");
           $stop; end
           end
  
       if(t==11) begin
           if(test_phase== 4'b1110)
           $display ("Output Verified");
           else begin
           $display ("Error");
           $stop; end
           end
 
       if(t==12) begin
           if(test_phase== 4'b1100)
           $display ("Output Verified");
           else begin
           $display ("Error");
           $stop; end
           end

       if(t==13) begin
           if(test_phase== 4'b1101)
           $display ("Output Verified");
           else begin
           $display ("Error"); 
           $stop; end
           end

       if(t==14) begin
           if(test_phase== 4'b1001)
           $display("Output Verified");
           else begin 
           $display ("Error");
           $stop; end
           end

       if(t==15) begin
           if(test_phase== 4'b1011)
           $display ("Output Verified");
           else begin
           $display ("Error");
           $stop; end
           end

       if(t==16) begin
           if(test_phase== 4'b0011)
           $display ("Output Verified");
           else begin 
           $display ("Error");
           $stop; end
           end

       if(t==17) begin
           if(test_phase== 4'b0111)
           $display ("Output Verified");
           else begin 
           $display ("Error"); 
           $stop; end
           end

       if(t==18) begin
           if(test_phase== 4'b0111)
           $display ("Output Verified");
           else begin
           $display ("Error"); 
           $stop; end
           end

       if(t==19) begin
           if(test_phase== 4'b0011)
           $display ("Output Verified");
           else begin 
           $display ("Error"); 
           $stop; end
           end

       if(t==20) begin
           if(test_phase== 4'b0011)
           $display ("Output Verified");
           else begin 
           $display ("Error");
           $stop; end
           end

       if(t==21) begin
           if(test_phase== 4'b1011)
           $display ("Output Verified");
           else begin 
           $display ("Error");
           $stop; end
           end

       if(t==22) begin
           if(test_phase== 4'b1011)
           $display ("Output Verified");
           else begin 
           $display ("Error");
           $stop; end
           end

       if(t==23) begin
           if(test_phase== 4'b1001)
           $display ("Output Verified");
           else begin
           $display ("Error"); 
           $stop; end
           end
                  
       if(t==24) begin
           if(test_phase== 4'b1001)
           $display ("Output Verified");
           else begin 
           $display ("Error"); 
           $stop; end
           end
                 
       if(t==25) begin
           if(test_phase== 4'b1101)
           $display ("Output Verified");
           else begin
           $display ("Error"); 
           $stop; end
           end
                 
       if(t==26) begin
           if(test_phase== 4'b1101)
           $display ("Output Verified");
           else begin 
           $display ("Error");
           $stop; end
           end            
                       
       if(t==27) begin
           if(test_phase== 4'b1100)
           $display ("Output Verified");
           else begin 
           $display ("Error");
           $stop; end
           end
               
       if(t==28) begin
           if(test_phase== 4'b1100)
           $display ("Output Verified");
           else begin 
           $display ("Error");
           $stop; end
           end
               
       if(t==29) begin
           if(test_phase== 4'b1110)
           $display ("Output Verified");
           else begin
           $display ("Error"); 
           $stop; end
           end
              
       if(t==30) begin
           if(test_phase== 4'b1110)
           $display ("Output Verified");
           else begin
           $display ("Error");
           $stop; end
           end
             
       if(t==31) begin
           if(test_phase== 4'b0110)
           $display ("Output Verified");
           else begin 
           $display ("Error");
           $stop; end
           end
                    
       if(t==32) begin
           if(test_phase== 4'b0110)
           $display ("Output Verified");
           else begin 
           $display ("Error");
           $stop; end
           end
                   
       if(t==33) begin
           if(test_phase== 4'b0111)
           $display ("Output Verified");
           else begin 
           $display ("Error");
           $stop; end
           end
           
       if(t==34) begin
           if(test_phase== 4'b0111)
           $display ("Output Verified");
           else begin 
           $display ("Error");
           $stop; end
           end
          
       if(t==35) begin
           if(test_phase== 4'b0011)
           $display ("Output Verified");
           else begin 
           $display ("Error"); 
           $stop; end
           end
         
       if(t==36) begin
           if(test_phase== 4'b0011)
           $display ("Output Verified");
           else begin 
           $display ("Error");
           $stop; end
           end
         
       if(t==37) begin
           if(test_phase== 4'b0111)
           $display ("Output Verified");
           else begin 
           $display ("Error");
           $stop; end
           end
       
       if(t==38) begin
           if(test_phase== 4'b0111)
           $display ("Output Verified");
           else begin
           $display ("Error");
           $stop; end
           end
       
       if(t==39) begin
           if(test_phase== 4'b0110)
           $display ("Output Verified");
           else begin 
           $display ("Error");
           $stop; end
           end 
     
       if(t==40) begin
           if(test_phase== 4'b0110)
           $display ("Output Verified");
           else begin 
           $display ("Error"); 
           $stop; end
           end
    
       if(t==41) begin
           if(test_phase== 4'b1110)
           $display ("Output Verified");
           else begin
           $display ("Error");
           $stop; end
           end
    
       if(t==42) begin
           if(test_phase== 4'b1110)
           $display ("Output Verified");
           else begin 
           $display ("Error");
           $stop; end
           end
     
       if(t==43) begin
           if(test_phase== 4'b1100)
           $display ("Output Verified");
           else begin 
           $display ("Error");
           $stop; end
           end
      
       if(t==44) begin
           if(test_phase== 4'b1100)
           $display ("Output Verified");
           else begin
           $display ("Error");
           $stop; end
           end
  
       if(t==45) begin
           if(test_phase== 4'b1101)
           $display ("Output Verified");
           else begin 
           $display ("Error");
           $stop; end
           end
   
       if(t==46) begin
           if(test_phase== 4'b1101)
           $display ("Output Verified");
           else begin 
           $display ("Error");
           $stop; end
           end 
     
       if(t==47) begin
           if(test_phase== 4'b1001)
           $display ("Output Verified");
           else begin 
           $display ("Error");
           $stop; end
           end
   
       if(t==48) begin
           if(test_phase== 4'b1001)
           $display ("Output Verified");
           else begin 
           $display ("Error"); 
           $stop; end
           end
   
       if(t==49) begin
           if(test_phase== 4'b1011)
           $display ("Output Verified");
           else begin 
           $display ("Error");
           $stop; end
           end
    
       if(t==50) begin
           if(test_phase== 4'b1011)
           $display ("Output Verified");
           else begin 
           $display ("Error");
           $stop; end                
           end
   
       if(t==51) begin
           if(test_phase== 4'b0011)
           $display ("Output Verified");
           else begin 
           $display ("Error");
           $stop; end 
           end

       if(t==52) begin
           if(test_phase== 4'b0011)
           $display ("Output Verified");
           else begin
           $display ("Error");
           $stop; end                
           end
   
       if(t==53) begin
           if(test_phase== 4'b0111)
           $display ("Output Verified");
           else begin 
           $display ("Error"); 
           $stop; end                    
           end
   
       if(t==54) begin
           if(test_phase== 4'b0111)
           begin
           $display ("Output Verified");
           $display ("ALL TESTS PASSED");
           end
           else begin 
           $display ("Error");
           $stop; end
           
           $stop;         
           end
 
       end  
   end      

endmodule
 
/********************************************************************************************************************
* Module ufmclk is the module which gets the clock from the oscillator
********************************************************************************************************************/

`timescale 1 ps / 1 ps                           
//synopsys translate_on
module  ufmclk_altufm_osc_7p3
	( 
	osc,
	oscena) /* synthesis synthesis_clearbox=1 */;
	output   osc;
	input   oscena;

	wire  wire_maxii_ufm_block1_osc;

	maxii_ufm   maxii_ufm_block1
	( 
	.arclk(1'b0),
	.ardin(1'b0),
	.arshft(1'b0),
	.bgpbusy(),
	.busy(),
	.drclk(1'b0),
	.drdout(),
	.drshft(1'b0),
	.osc(wire_maxii_ufm_block1_osc),
	.oscena(oscena)
	`ifdef FORMAL_VERIFICATION
	`else
	// synopsys translate_off
	`endif
	,
	.drdin(1'b0),
	.erase(1'b0),
	.program(1'b0)
	`ifdef FORMAL_VERIFICATION
	`else
	// synopsys translate_on
	`endif
	// synopsys translate_off
	,
	.ctrl_bgpbusy(),
	.devclrn(),
	.devpor(),
	.sbdin(),
	.sbdout()
	// synopsys translate_on
	);
	defparam
		maxii_ufm_block1.address_width = 9,
		maxii_ufm_block1.osc_sim_setting = 180000,
		maxii_ufm_block1.lpm_type = "maxii_ufm";
	assign
		osc = wire_maxii_ufm_block1_osc;
endmodule //ufmclk_altufm_osc_7p3
//VALID FILE


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module ufmclk (
	oscena,
	osc)/* synthsim:/testbench/t
esis synthesis_clearbox = 1 */;

	input	  oscena;
	output	  osc;

	wire  sub_wire0;
	wire  osc = sub_wire0;

	ufmclk_altufm_osc_7p3	ufmclk_altufm_osc_7p3_component (
				.oscena (oscena),
				.osc (sub_wire0));

endmodule

/***************************************************************************************************************************
* module divider divides the clock from ufmclk to produce a 
  clock suitable to drive the motor controller 
***************************************************************************************************************************/
 module divider1 (osc, clk,clk1);                 
	   input osc;
   	   output clk,clk1;
   	   reg clk,clk1;
       reg [16:0] count;
 initial
       count= 17'b00000000000000000;

 always @( posedge osc)
      begin
         count = count + 1;
         clk = count[16];
         clk1=count[15];
      end

endmodule

/********************************** END ********************************************************************************/
