library verilog;
use verilog.vl_types.all;
entity ufmclk_altufm_osc_7p3 is
    port(
        osc             : out    vl_logic;
        oscena          : in     vl_logic
    );
end ufmclk_altufm_osc_7p3;
