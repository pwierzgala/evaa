library verilog;
use verilog.vl_types.all;
entity MAXII_PRIM_DFFE is
    // This module cannot be connected to from
    // VHDL because it has unnamed ports.
end MAXII_PRIM_DFFE;
